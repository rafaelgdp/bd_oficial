module AMBA(
	input logic valid,
	input logic [7:0] data_in,
	input logic [7:0] address,
	output logic [7:0] data_out,
	output logic ready
);



endmodule
