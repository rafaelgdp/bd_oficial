module RegisterField(
	input logic [7:0] DATA_0_IN,
	input logic [7:0] DATA_1_IN,
	input logic [7:0] ADDRESS,
	output logic [7:0] BD_DATA_0,
	output logic [7:0] BD_DATA_1
);

logic [7:0] BD_CONTROL;
/*logic [7:0] BD_DATA_0;
logic [7:0] BD_DATA_1;*/

/*case address
x: bd_data_0 <= data; 
y: bd_data_1 <= data;*/

endmodule

