module RegisterField(
	input logic [7:0] DATA,
	input logic [7:0] ADDRESS
);

logic [7:0] BD_CONTROL;
logic [7:0] BD_DATA_0;
logic [7:0] BD_DATA_1;

endmodule

